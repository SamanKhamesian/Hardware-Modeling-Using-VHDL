LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY FIFO IS

	PORT(
	
		In_Data:	IN	STD_LOGIC_VECTOR(15 DOWNTO 0);
		Out_Data:	OUT	STD_LOGIC_VECTOR(15 DOWNTO 0);
		RST:		IN	STD_LOGIC;
		CLK:		IN	STD_LOGIC;
		EN:			IN	STD_LOGIC
	);
	
END FIFO;

ARCHITECTURE ARCH_FIFO OF FIFO IS
	
	SIGNAL	OUTPUT:		STD_LOGIC_VECTOR(15 DOWNTO 0);
	TYPE	MEM_TYPE 	IS ARRAY(0 TO 3) OF STD_LOGIC_VECTOR(15 DOWNTO 0);
	SIGNAL	FIFO_MEM:	MEM_TYPE:= (OTHERS => (OTHERS => '0'));
	
BEGIN
	
	PROCESS (CLK, RST) BEGIN
	
		IF (RST = '1') THEN
		
			OUTPUT		<= (OTHERS => '0');
			FIFO_MEM	<= (OTHERS => (OTHERS => '0'));

		ELSIF (RISING_EDGE(CLK) AND EN = '1') THEN
		
			OUTPUT		<= FIFO_MEM(3);
			FIFO_MEM(3)	<= FIFO_MEM(2);
			FIFO_MEM(2) <= FIFO_MEM(1);
			FIFO_MEM(1) <= FIFO_MEM(0);
			FIFO_MEM(0) <= In_Data;
				
		END IF;
			
	END PROCESS;
	
	Out_Data <= OUTPUT;

END ARCH_FIFO;
